`define NOP 3'b000
`define ADD 3'b010
`define ADDI 3'b110
`define MULI 3'b111
`define LOAD 3'b100
