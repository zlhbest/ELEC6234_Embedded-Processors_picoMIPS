`define RI 2'b00
`define ADD 2'b10
`define MUL 2'b11
